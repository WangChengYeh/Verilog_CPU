// 指令編碼
`define OPCODE_LOAD    3'b000
`define OPCODE_STORE   3'b001
`define OPCODE_ADD     3'b010
`define OPCODE_CMP     3'b011
`define OPCODE_JUMP    3'b100